module top ();


A module A();
B module B();

//module A();
//Critical path Logic()

//module B();
//Non critical path logic()
endmodule