module top ();

Critical path Logic()
Non critical path logic()
endmodule